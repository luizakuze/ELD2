--=============================
-- Listing 8.15 programmable mod-m counter
--=============================
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
entity prog_counter is
   port(
      clk, reset: in std_logic;
		clk_out: out std_logic;
      m: in std_logic_vector(3 downto 0);
      q: out std_logic_vector(3 downto 0)
   );
end prog_counter;

architecture two_seg_clear_arch of prog_counter is
   signal r_reg: unsigned(3 downto 0);
   signal r_next: unsigned(3 downto 0);
begin
   -- register
   process(clk,reset)
   begin
      if (reset='1') then
         r_reg <= (others=>'0');
      elsif (clk'event and clk='1') then
         r_reg <= r_next;
      end if;
   end process;
   -- next-state logic
   r_next <= (others=>'0') when r_reg=(unsigned(m)-1) else
             r_reg + 1;
   -- output logic
   q <= std_logic_vector(r_reg);
	clk_out <= '1' when r_reg=((unsigned(m)-1)/2) else '0';
end two_seg_clear_arch;


--=============================
-- Listing 8.16
--=============================
architecture two_seg_effi_arch of prog_counter is
   signal r_reg: unsigned(3 downto 0);
   signal r_next, r_inc: unsigned(3 downto 0);
begin
   -- register
   process(clk,reset)
   begin
      if (reset='1') then
         r_reg <= (others=>'0');
      elsif (clk'event and clk='1') then
         r_reg <= r_next;
      end if;
   end process;
   -- next-state logic
   r_inc <= r_reg + 1;
   r_next <= (others=>'0') when r_inc=unsigned(m) else
             r_inc;
   -- output logic
   q <= std_logic_vector(r_reg);
end two_seg_effi_arch;


configuration cfg_ifsc of prog_counter is  
	for two_seg_clear_arch end for;
--for two_seg_effi_arch end for;
end cfg_ifsc;
